//20L152 SUMITHA R A

module halfadd(
    input a,b,
    output s,co
    );
assign s=a^b;
assign co=a&b;

endmodule


